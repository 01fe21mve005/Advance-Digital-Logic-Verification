//class monitor

class monitor

int no_repeat count;
mail box mon2scb;

function(mailbox mon2scd)
this.mon2scb=mon2scb;
endfunction

task main()


if(trans data 

