//interface.sv

class interface

logic bit [1:0] data;
logic bit [1:0] addr;
logic bit [1:0] addr a;
logic bit [1:0] addr b;
logic bit [1:0] data a;
logic bit [1:0] data b;

end class 
